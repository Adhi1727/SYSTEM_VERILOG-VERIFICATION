# KERNEL: ASDB file was created in location /home/runner/dataset.asdb
# KERNEL: GENERATOR CHECKED
# KERNEL:                    0rst = 0 | d = 1 | q = 0
# KERNEL: DRIVER CHECKED
# KERNEL:                    5rst = 0 | d = 1 | q = 0
# KERNEL: rst = 1
# KERNEL: MONITOR CHECKED
# KERNEL:                    5rst = 1 | d = 0 | q = 0
# KERNEL: SCOREBOARD CHECKED
# KERNEL:                    5rst = 1 | d = 0 | q = 0
# KERNEL: Result : pass
# KERNEL: GENERATOR CHECKED
# KERNEL:                    5rst = 0 | d = 1 | q = 0
# KERNEL: MONITOR CHECKED
# KERNEL:                   15rst = 1 | d = 1 | q = 0
# KERNEL: DRIVER CHECKED
# KERNEL:                   15rst = 0 | d = 1 | q = 0
# KERNEL: rst = 1
# KERNEL: SCOREBOARD CHECKED
# KERNEL:                   15rst = 1 | d = 1 | q = 0
# KERNEL: Result : pass
# KERNEL: GENERATOR CHECKED
# KERNEL:                   15rst = 0 | d = 0 | q = 0
# KERNEL: MONITOR CHECKED
# KERNEL:                   25rst = 0 | d = 1 | q = 1
# KERNEL: DRIVER CHECKED
# KERNEL:                   25rst = 0 | d = 0 | q = 0
# KERNEL: rst = 0
# KERNEL: SCOREBOARD CHECKED
# KERNEL:                   25rst = 0 | d = 1 | q = 1
# KERNEL: Result : pass
# KERNEL: GENERATOR CHECKED
# KERNEL:                   25rst = 0 | d = 1 | q = 0
# KERNEL: MONITOR CHECKED
# KERNEL:                   35rst = 0 | d = 0 | q = 0
# KERNEL: DRIVER CHECKED
# KERNEL:                   35rst = 0 | d = 1 | q = 0
# KERNEL: rst = 0
# KERNEL: SCOREBOARD CHECKED
# KERNEL:                   35rst = 0 | d = 0 | q = 0
# KERNEL: Result : pass
# KERNEL: GENERATOR CHECKED
# KERNEL:                   35rst = 0 | d = 1 | q = 0
# KERNEL: MONITOR CHECKED
# KERNEL:                   45rst = 0 | d = 1 | q = 1
# KERNEL: DRIVER CHECKED
# KERNEL:                   45rst = 0 | d = 1 | q = 0
# KERNEL: rst = 0
# KERNEL: SCOREBOARD CHECKED
# KERNEL:                   45rst = 0 | d = 1 | q = 1
# KERNEL: Result : pass
# RUNTIME: Info: RUNTIME_0068 $finish called.
