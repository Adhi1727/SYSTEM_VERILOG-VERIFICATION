interface inter;
  logic clk;
  logic r_w;
  logic [3:0]addr;
  logic [7:0]wr_d;
  logic [7:0]rd_d;
endinterface
